module tst();
endmodule
module tst2();
endmodule
module tst3();
endmodule
