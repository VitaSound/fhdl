`include "foo.v"
`include "bar.v"
`include "baz.v"
module tst1(a, b, c);
endmodule
module tst2();
endmodule
module tst3();
endmodule
