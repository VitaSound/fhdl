module tst1;
a port,
b port,
a port,

endmodule
module tst2;

endmodule
