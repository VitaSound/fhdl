module tst
endmodule
